--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:38:39 10/21/2019
-- Design Name:   
-- Module Name:   C:/Users/Dell/Documents/aprender vhdl/contadorcomonolivro/contadorcomonolivro_tb.vhd
-- Project Name:  contadorcomonolivro
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: contadorsimples
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY contadorcomonolivro_tb IS
END contadorcomonolivro_tb;
 
ARCHITECTURE behavior OF contadorcomonolivro_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT contadorsimples
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         ena : IN  std_logic;
         full_count : OUT  std_logic;
         dig1 : OUT  std_logic_vector(6 downto 0);
         dig2 : OUT  std_logic_vector(6 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal ena : std_logic := '0';

 	--Outputs
   signal full_count : std_logic;
   signal dig1 : std_logic_vector(6 downto 0);
   signal dig2 : std_logic_vector(6 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: contadorsimples PORT MAP (
          clk => clk,
          rst => rst,
          ena => ena,
          full_count => full_count,
          dig1 => dig1,
          dig2 => dig2
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
      ena<='1';
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
