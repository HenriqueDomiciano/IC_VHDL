
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:38:23 09/03/2019 
-- Design Name: 
-- Module Name:    testadordeprioridade - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testadordeprioridade is
port( a : in std_logic_vector (7 downto 0);
		b : out std_logic_vector (7 downto 0)
);
end testadordeprioridade;

architecture Behavioral of testadordeprioridade is
begin

when a(7)='1' 
end Behavioral;

