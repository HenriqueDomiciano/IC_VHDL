--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package packageforarray is
type matrix is array (natural range<>,natural range <>) of std_logic;
end packageforarray;

package body packageforarray is
 end packageforarray;
