----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:23:02 09/30/2019 
-- Design Name: 
-- Module Name:    registradordedeslocamento - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity registradordedeslocamento is
	port(
													)
end registradordedeslocamento;

architecture Behavioral of registradordedeslocamento is

begin


end Behavioral;

